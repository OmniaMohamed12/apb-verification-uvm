package APB_Pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "APB_Sequence_Item.svh"
    `include "APB_SequenceS.svh"
    `include "APB_Sequencer.svh"
    `include "APB_Driver.svh"
    `include "APB_Monitor.svh"
    `include "APB_Agent.svh"
    `include "APB_Scoreboard.svh"
    `include "APB_Coverage.svh"
    `include "APB_Env.svh"
    `include "APB_Test.svh"

endpackage